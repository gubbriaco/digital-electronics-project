library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package MyDefinitions is

    constant n: integer:=16; -- numero di bit da sommare
    constant nFA: integer:= n/2; -- numero di Full-Adder per blocco

end package;
