library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package MyDefinitions is
    constant n_bit: integer:=16;
end package;